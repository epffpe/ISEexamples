--
-- Definition of a single port ROM for KCPSM3 program defined by monitor.psm
-- and assmbled using KCPSM3 assembler.
--
-- Standard IEEE libraries
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
--
-- The Unisim Library is used to define Xilinx primitives. It is also used during
-- simulation. The source can be viewed at %XILINX%\vhdl\src\unisims\unisim_VCOMP.vhd
--  
library unisim;
use unisim.vcomponents.all;
--
--
entity monitor is
    Port (      address : in std_logic_vector(9 downto 0);
            instruction : out std_logic_vector(17 downto 0);
                    clk : in std_logic);
    end monitor;
--
architecture low_level_definition of monitor is
--
-- Attributes to define ROM contents during implementation synthesis. 
-- The information is repeated in the generic map for functional simulation
--
attribute INIT_00 : string; 
attribute INIT_01 : string; 
attribute INIT_02 : string; 
attribute INIT_03 : string; 
attribute INIT_04 : string; 
attribute INIT_05 : string; 
attribute INIT_06 : string; 
attribute INIT_07 : string; 
attribute INIT_08 : string; 
attribute INIT_09 : string; 
attribute INIT_0A : string; 
attribute INIT_0B : string; 
attribute INIT_0C : string; 
attribute INIT_0D : string; 
attribute INIT_0E : string; 
attribute INIT_0F : string; 
attribute INIT_10 : string; 
attribute INIT_11 : string; 
attribute INIT_12 : string; 
attribute INIT_13 : string; 
attribute INIT_14 : string; 
attribute INIT_15 : string; 
attribute INIT_16 : string; 
attribute INIT_17 : string; 
attribute INIT_18 : string; 
attribute INIT_19 : string; 
attribute INIT_1A : string; 
attribute INIT_1B : string; 
attribute INIT_1C : string; 
attribute INIT_1D : string; 
attribute INIT_1E : string; 
attribute INIT_1F : string; 
attribute INIT_20 : string; 
attribute INIT_21 : string; 
attribute INIT_22 : string; 
attribute INIT_23 : string; 
attribute INIT_24 : string; 
attribute INIT_25 : string; 
attribute INIT_26 : string; 
attribute INIT_27 : string; 
attribute INIT_28 : string; 
attribute INIT_29 : string; 
attribute INIT_2A : string; 
attribute INIT_2B : string; 
attribute INIT_2C : string; 
attribute INIT_2D : string; 
attribute INIT_2E : string; 
attribute INIT_2F : string; 
attribute INIT_30 : string; 
attribute INIT_31 : string; 
attribute INIT_32 : string; 
attribute INIT_33 : string; 
attribute INIT_34 : string; 
attribute INIT_35 : string; 
attribute INIT_36 : string; 
attribute INIT_37 : string; 
attribute INIT_38 : string; 
attribute INIT_39 : string; 
attribute INIT_3A : string; 
attribute INIT_3B : string; 
attribute INIT_3C : string; 
attribute INIT_3D : string; 
attribute INIT_3E : string; 
attribute INIT_3F : string; 
attribute INITP_00 : string;
attribute INITP_01 : string;
attribute INITP_02 : string;
attribute INITP_03 : string;
attribute INITP_04 : string;
attribute INITP_05 : string;
attribute INITP_06 : string;
attribute INITP_07 : string;
--
-- Attributes to define ROM contents during implementation synthesis.
--
attribute INIT_00 of ram_1024_x_18  : label is "E00CE00BE00AE009E008E007E006E005E004E003E002E001E0000000C08000FF";
attribute INIT_01 of ram_1024_x_18  : label is "4041509E40545017400D01BE013001EC0259C0010C000D00E006000C0167E00D";
attribute INIT_02 of ram_1024_x_18  : label is "007A40170231502F405750614052517A4050512340425145405350EC404C50B7";
attribute INIT_03 of ram_1024_x_18  : label is "130001BE1600585B03D8120001BE130001BE542D402001BE58770088505E4A00";
attribute INIT_04 of ram_1024_x_18  : label is "C980E980C980E980C660C980F9A009ED542D400D01BE1500585B03D8120001BE";
attribute INIT_05 of ram_1024_x_18  : label is "028F02694017028602694017C98000FFC980E980C980E980C560C980F9A009F6";
attribute INIT_06 of ram_1024_x_18  : label is "F9A009B603C14004C980F9A009AD542D400D01BE58770088505E4A00007A4017";
attribute INIT_07 of ram_1024_x_18  : label is "B400402001BE120001BE0A004017027902694017020DC98000FF03C14004C980";
attribute INIT_08 of ram_1024_x_18  : label is "01BEC014B800D2000203B80003E501BEA0000A20A0000A04B400424250864241";
attribute INIT_09 of ram_1024_x_18  : label is "404901BEA000C011B80003D8120001BE130001BEC012B80003D8120001BE1300";
attribute INIT_0A of ram_1024_x_18  : label is "5817019B542D4020401701D154AC400D01BE542D404501BE542D404D01BE542D";
attribute INIT_0B of ram_1024_x_18  : label is "542D405201BE542D404101BE542D404C01BE401701D1E005E004E408E507E606";
attribute INIT_0C of ram_1024_x_18  : label is "5817019BC10150D5404F01BE542D4020401701D554C8400D01BE542D404D01BE";
attribute INIT_0D of ram_1024_x_18  : label is "401701D5E00CC002600C542D400D01BE54E0404E01BE401701D5E40BE50AE609";
attribute INIT_0E of ram_1024_x_18  : label is "01BE542D404501BE401701D5E00C0000542D400D01BE542D404601BE542D4046";
attribute INIT_0F of ram_1024_x_18  : label is "40FC0A065900C0010A015D1F8008591F80C84017016A54F7400D01BE542D4044";
attribute INIT_10 of ram_1024_x_18  : label is "0167E00DD0A0600D542D400D01BE5511404E01BE542D404F01BE542D402001BE";
attribute INIT_11 of ram_1024_x_18  : label is "026940170167E00DB0A0EAFF600D542D400D01BE542D404601BE542D40464017";
attribute INIT_12 of ram_1024_x_18  : label is "01BE542D404F01BE542D405401BE542D405401BE542D405501BE4017020D02DB";
attribute INIT_13 of ram_1024_x_18  : label is "414102AA59400A0C021001CA8F301FB002CF0B004A03542D400D01BE542D404E";
attribute INIT_14 of ram_1024_x_18  : label is "404301BE542D405401BE542D404901BE542D405701BE401755374B048B0102B0";
attribute INIT_15 of ram_1024_x_18  : label is "59620A0C021001CA8F301FB002C20B004A02542D400D01BE542D404801BE542D";
attribute INIT_16 of ram_1024_x_18  : label is "01CA8F301FB002DB0B006A0DA000C0A0600D401755594B088B0102B0416302AA";
attribute INIT_17 of ram_1024_x_18  : label is "542D404F01BE542D405201BEA000556C4B088B0102B0417602AA59750A0C0210";
attribute INIT_18 of ram_1024_x_18  : label is "5999EB00CA010AFF0BFFC0400000C0400001020D542D400D01BE542D404D01BE";
attribute INIT_19 of ram_1024_x_18  : label is "01BE8101162059B903B340170216418B01CA519A4FFF4F05518D202040000307";
attribute INIT_1A of ram_1024_x_18  : label is "55B9400D01BE8101142059B903B355B9403A01BE8101152059B903B355B9403A";
attribute INIT_1B of ram_1024_x_18  : label is "03A97010A000000E000102960269A000000E00005DB9443C5DB9453C5DB94618";
attribute INIT_1C of ram_1024_x_18  : label is "CFC041CA030751CF20024000A00001CA4F0141C2030755C720104000A0008101";
attribute INIT_1D of ram_1024_x_18  : label is "2002A00002B551DF2001600C0210029F01E502E20E09A00001E502E20E06A000";
attribute INIT_1E of ram_1024_x_18  : label is "400082101210013041E68101B0004F0D01CA7F100130A00002AAA00002B051E3";
attribute INIT_1F of ram_1024_x_18  : label is "02105A024130C101021355EF5120810151FC4F08B0004F0DFF1001C256042008";
attribute INIT_20 of ram_1024_x_18  : label is "A00001CA0F0D42084F01B00020104000020D023EEF30020D41EC026641EF0213";
attribute INIT_21 of ram_1024_x_18  : label is "01CA0F6B01CA0F6301CA0F6501CA0F6801CA0F43A00001CA0F08A00001CA0F20";
attribute INIT_22 of ram_1024_x_18  : label is "01CA0F6B01CA0F6E01CA0F6901CA0F6C021001CA0F3101CA0F5001CA0F4A0210";
attribute INIT_23 of ram_1024_x_18  : label is "01CA0F4F424E01CA0F7801CA0F6101CA0F7401CA0F6E01CA0F7901CA0F53420D";
attribute INIT_24 of ram_1024_x_18  : label is "0F45021001CA0F7701CA0F6F01CA0F6C01CA0F6601CA0F7201CA0F6501CA0F76";
attribute INIT_25 of ram_1024_x_18  : label is "01CA0F5001CA0F4301CA0F4B020D420D01CA0F7201CA0F6F01CA01CA0F7201CA";
attribute INIT_26 of ram_1024_x_18  : label is "0F6101CA0F7601CA0F6E01CA0F49A00001CA0F3E01CA0F3301CA0F4D01CA0F53";
attribute INIT_27 of ram_1024_x_18  : label is "01CA0F7201CA01CA0F6401CA0F41A000021001CA0F6401CA0F6901CA0F6C01CA";
attribute INIT_28 of ram_1024_x_18  : label is "0F52420D01CA0F6101CA0F7401CA0F6101CA0F44420D01CA01CA0F7301CA0F65";
attribute INIT_29 of ram_1024_x_18  : label is "0F41420D01CA0F6501CA0F6D01CA0F6901CA0F54420D01CA0F4D01CA0F4101CA";
attribute INIT_2A of ram_1024_x_18  : label is "420D01CA01CA0F4601CA0F4FA00001CA0F6D01CA0F7201CA0F6101CA0F6C01CA";
attribute INIT_2B of ram_1024_x_18  : label is "0F6501CA0F7601CA0F6901CA0F7401CA0F6301CA0F41420D01CA0F4E01CA0F4F";
attribute INIT_2C of ram_1024_x_18  : label is "0F42A00001CA0F6801CA0F6301CA0F7401CA0F6901CA0F7701CA0F53420D01CA";
attribute INIT_2D of ram_1024_x_18  : label is "0F4401CA0F4501CA0F4CA00001CA0F6E01CA0F6F01CA01CA0F7401CA0F7501CA";
attribute INIT_2E of ram_1024_x_18  : label is "F120030070E08E018201F020003A8201F0208201F120030070E00230A00001CA";
attribute INIT_2F of ram_1024_x_18  : label is "A000F020000D8201F0208201F120030070E08E018201F020003A8201F0208201";
attribute INIT_30 of ram_1024_x_18  : label is "C00063016200E515E414E313E212E111E010A000803AC1015F01C00A81010130";
attribute INIT_31 of ram_1024_x_18  : label is "80015B21E303C2E80000B350924063036202F530D42065016400C001EC01ED00";
attribute INIT_32 of ram_1024_x_18  : label is "82E8433180015B2FE303C2E80000A300920063056204E303E202A30382E8431C";
attribute INIT_33 of ram_1024_x_18  : label is "E1075341413C81016107E1080100434BE1085339413C91006108E305E204A303";
attribute INIT_34 of ram_1024_x_18  : label is "6007575C501061096006E1060100434BE1065349411881016106E1070100434B";
attribute INIT_35 of ram_1024_x_18  : label is "53612001600C05FFE00CC001535C2002600C575C5010610B6008575C5010610A";
attribute INIT_36 of ram_1024_x_18  : label is "C2E2B2400389800AC1015F68C00A810101006006047F53662002600504FF057F";
attribute INIT_37 of ram_1024_x_18  : label is "03891010C2E0B2500389800AC1015F76C00A810101006007C2E3B25003891010";
attribute INIT_38 of ram_1024_x_18  : label is "02A4B800C00102F9B800C00102C0A000651564146313621261116010C2E1B250";
attribute INIT_39 of ram_1024_x_18  : label is "C00102F8B800C0010282B800C0010292B800C0010299B800C00102B0B800C001";
attribute INIT_3A of ram_1024_x_18  : label is "80C6A000A0DFBC00407BB8004061A00002FFB800C0010290B800C0010280B800";
attribute INIT_3B of ram_1024_x_18  : label is "9200B80003AF7010810102069200020602061200B80003AF7010A000C0F6B800";
attribute INIT_3C of ram_1024_x_18  : label is "A00F1010120003D3000E000E000E000E1100A00001CA1F1001CA1F2003C7A000";
attribute INIT_3D of ram_1024_x_18  : label is "03060306030603061300B80003E51030A000803A80075BD6C00AA000110003D3";
attribute INIT_3E of ram_1024_x_18  : label is "800AA000C0F6B80080075FEFC011B800C0E9B80080B9A000D030B80003E51020";
attribute INIT_3F of ram_1024_x_18  : label is "43FC8001AC008D0100000000000000000000000000000000000000000000A000";
attribute INITP_00 of ram_1024_x_18 : label is "9CCFFE320C837FDFFFF888A088A0DCF333CCF7FDFF7777777773F08EAAAAAA88";
attribute INITP_01 of ram_1024_x_18 : label is "ED377F7DF7F8DF7DF837DFEAF77DFDF7DF7DFEAAFDFDF7DF7AB33ACCE92F889D";
attribute INITP_02 of ram_1024_x_18 : label is "DF7B5FFBD30A3D7FEF4C37DF7DF7DFD7FEF4C37DF7DF7DFFFE037DF7E0DF7DF7";
attribute INITP_03 of ram_1024_x_18 : label is "F5F5D9BD10D9C2EF6F4FF2F2BF4B3F49CA3E8DDDDD3F74FDD3FFF4D3D4223DF7";
attribute INITP_04 of ram_1024_x_18 : label is "CF32F3333332CCCCCCCFCCF33CCCCCCCCF333333CCCCF333CCCCCB2CB324FBFF";
attribute INITP_05 of ram_1024_x_18 : label is "A19B1619B1619B0B332CCF332CCCCCCF333333CCFCCB33333CCCCF333CCCCFCC";
attribute INITP_06 of ram_1024_x_18 : label is "C8D7508C8D750340D08D34343423B523B523B529775142977514143AC2AAA5D4";
attribute INITP_07 of ram_1024_x_18 : label is "F50000026676662CAA2C976303AA2CCE6C668B26626624924924924924920008";
--
begin
--
  --Instantiate the Xilinx primitive for a block RAM
  ram_1024_x_18: RAMB16_S18
  --synthesis translate_off
  --INIT values repeated to define contents for functional simulation
  generic map ( INIT_00 => X"E00CE00BE00AE009E008E007E006E005E004E003E002E001E0000000C08000FF",
                INIT_01 => X"4041509E40545017400D01BE013001EC0259C0010C000D00E006000C0167E00D",
                INIT_02 => X"007A40170231502F405750614052517A4050512340425145405350EC404C50B7",
                INIT_03 => X"130001BE1600585B03D8120001BE130001BE542D402001BE58770088505E4A00",
                INIT_04 => X"C980E980C980E980C660C980F9A009ED542D400D01BE1500585B03D8120001BE",
                INIT_05 => X"028F02694017028602694017C98000FFC980E980C980E980C560C980F9A009F6",
                INIT_06 => X"F9A009B603C14004C980F9A009AD542D400D01BE58770088505E4A00007A4017",
                INIT_07 => X"B400402001BE120001BE0A004017027902694017020DC98000FF03C14004C980",
                INIT_08 => X"01BEC014B800D2000203B80003E501BEA0000A20A0000A04B400424250864241",
                INIT_09 => X"404901BEA000C011B80003D8120001BE130001BEC012B80003D8120001BE1300",
                INIT_0A => X"5817019B542D4020401701D154AC400D01BE542D404501BE542D404D01BE542D",
                INIT_0B => X"542D405201BE542D404101BE542D404C01BE401701D1E005E004E408E507E606",
                INIT_0C => X"5817019BC10150D5404F01BE542D4020401701D554C8400D01BE542D404D01BE",
                INIT_0D => X"401701D5E00CC002600C542D400D01BE54E0404E01BE401701D5E40BE50AE609",
                INIT_0E => X"01BE542D404501BE401701D5E00C0000542D400D01BE542D404601BE542D4046",
                INIT_0F => X"40FC0A065900C0010A015D1F8008591F80C84017016A54F7400D01BE542D4044",
                INIT_10 => X"0167E00DD0A0600D542D400D01BE5511404E01BE542D404F01BE542D402001BE",
                INIT_11 => X"026940170167E00DB0A0EAFF600D542D400D01BE542D404601BE542D40464017",
                INIT_12 => X"01BE542D404F01BE542D405401BE542D405401BE542D405501BE4017020D02DB",
                INIT_13 => X"414102AA59400A0C021001CA8F301FB002CF0B004A03542D400D01BE542D404E",
                INIT_14 => X"404301BE542D405401BE542D404901BE542D405701BE401755374B048B0102B0",
                INIT_15 => X"59620A0C021001CA8F301FB002C20B004A02542D400D01BE542D404801BE542D",
                INIT_16 => X"01CA8F301FB002DB0B006A0DA000C0A0600D401755594B088B0102B0416302AA",
                INIT_17 => X"542D404F01BE542D405201BEA000556C4B088B0102B0417602AA59750A0C0210",
                INIT_18 => X"5999EB00CA010AFF0BFFC0400000C0400001020D542D400D01BE542D404D01BE",
                INIT_19 => X"01BE8101162059B903B340170216418B01CA519A4FFF4F05518D202040000307",
                INIT_1A => X"55B9400D01BE8101142059B903B355B9403A01BE8101152059B903B355B9403A",
                INIT_1B => X"03A97010A000000E000102960269A000000E00005DB9443C5DB9453C5DB94618",
                INIT_1C => X"CFC041CA030751CF20024000A00001CA4F0141C2030755C720104000A0008101",
                INIT_1D => X"2002A00002B551DF2001600C0210029F01E502E20E09A00001E502E20E06A000",
                INIT_1E => X"400082101210013041E68101B0004F0D01CA7F100130A00002AAA00002B051E3",
                INIT_1F => X"02105A024130C101021355EF5120810151FC4F08B0004F0DFF1001C256042008",
                INIT_20 => X"A00001CA0F0D42084F01B00020104000020D023EEF30020D41EC026641EF0213",
                INIT_21 => X"01CA0F6B01CA0F6301CA0F6501CA0F6801CA0F43A00001CA0F08A00001CA0F20",
                INIT_22 => X"01CA0F6B01CA0F6E01CA0F6901CA0F6C021001CA0F3101CA0F5001CA0F4A0210",
                INIT_23 => X"01CA0F4F424E01CA0F7801CA0F6101CA0F7401CA0F6E01CA0F7901CA0F53420D",
                INIT_24 => X"0F45021001CA0F7701CA0F6F01CA0F6C01CA0F6601CA0F7201CA0F6501CA0F76",
                INIT_25 => X"01CA0F5001CA0F4301CA0F4B020D420D01CA0F7201CA0F6F01CA01CA0F7201CA",
                INIT_26 => X"0F6101CA0F7601CA0F6E01CA0F49A00001CA0F3E01CA0F3301CA0F4D01CA0F53",
                INIT_27 => X"01CA0F7201CA01CA0F6401CA0F41A000021001CA0F6401CA0F6901CA0F6C01CA",
                INIT_28 => X"0F52420D01CA0F6101CA0F7401CA0F6101CA0F44420D01CA01CA0F7301CA0F65",
                INIT_29 => X"0F41420D01CA0F6501CA0F6D01CA0F6901CA0F54420D01CA0F4D01CA0F4101CA",
                INIT_2A => X"420D01CA01CA0F4601CA0F4FA00001CA0F6D01CA0F7201CA0F6101CA0F6C01CA",
                INIT_2B => X"0F6501CA0F7601CA0F6901CA0F7401CA0F6301CA0F41420D01CA0F4E01CA0F4F",
                INIT_2C => X"0F42A00001CA0F6801CA0F6301CA0F7401CA0F6901CA0F7701CA0F53420D01CA",
                INIT_2D => X"0F4401CA0F4501CA0F4CA00001CA0F6E01CA0F6F01CA01CA0F7401CA0F7501CA",
                INIT_2E => X"F120030070E08E018201F020003A8201F0208201F120030070E00230A00001CA",
                INIT_2F => X"A000F020000D8201F0208201F120030070E08E018201F020003A8201F0208201",
                INIT_30 => X"C00063016200E515E414E313E212E111E010A000803AC1015F01C00A81010130",
                INIT_31 => X"80015B21E303C2E80000B350924063036202F530D42065016400C001EC01ED00",
                INIT_32 => X"82E8433180015B2FE303C2E80000A300920063056204E303E202A30382E8431C",
                INIT_33 => X"E1075341413C81016107E1080100434BE1085339413C91006108E305E204A303",
                INIT_34 => X"6007575C501061096006E1060100434BE1065349411881016106E1070100434B",
                INIT_35 => X"53612001600C05FFE00CC001535C2002600C575C5010610B6008575C5010610A",
                INIT_36 => X"C2E2B2400389800AC1015F68C00A810101006006047F53662002600504FF057F",
                INIT_37 => X"03891010C2E0B2500389800AC1015F76C00A810101006007C2E3B25003891010",
                INIT_38 => X"02A4B800C00102F9B800C00102C0A000651564146313621261116010C2E1B250",
                INIT_39 => X"C00102F8B800C0010282B800C0010292B800C0010299B800C00102B0B800C001",
                INIT_3A => X"80C6A000A0DFBC00407BB8004061A00002FFB800C0010290B800C0010280B800",
                INIT_3B => X"9200B80003AF7010810102069200020602061200B80003AF7010A000C0F6B800",
                INIT_3C => X"A00F1010120003D3000E000E000E000E1100A00001CA1F1001CA1F2003C7A000",
                INIT_3D => X"03060306030603061300B80003E51030A000803A80075BD6C00AA000110003D3",
                INIT_3E => X"800AA000C0F6B80080075FEFC011B800C0E9B80080B9A000D030B80003E51020",
                INIT_3F => X"43FC8001AC008D0100000000000000000000000000000000000000000000A000",    
               INITP_00 => X"9CCFFE320C837FDFFFF888A088A0DCF333CCF7FDFF7777777773F08EAAAAAA88",
               INITP_01 => X"ED377F7DF7F8DF7DF837DFEAF77DFDF7DF7DFEAAFDFDF7DF7AB33ACCE92F889D",
               INITP_02 => X"DF7B5FFBD30A3D7FEF4C37DF7DF7DFD7FEF4C37DF7DF7DFFFE037DF7E0DF7DF7",
               INITP_03 => X"F5F5D9BD10D9C2EF6F4FF2F2BF4B3F49CA3E8DDDDD3F74FDD3FFF4D3D4223DF7",
               INITP_04 => X"CF32F3333332CCCCCCCFCCF33CCCCCCCCF333333CCCCF333CCCCCB2CB324FBFF",
               INITP_05 => X"A19B1619B1619B0B332CCF332CCCCCCF333333CCFCCB33333CCCCF333CCCCFCC",
               INITP_06 => X"C8D7508C8D750340D08D34343423B523B523B529775142977514143AC2AAA5D4",
               INITP_07 => X"F50000026676662CAA2C976303AA2CCE6C668B26626624924924924924920008")
  --synthesis translate_on
  port map(    DI => "0000000000000000",
              DIP => "00",
               EN => '1',
               WE => '0',
              SSR => '0',
              CLK => clk,
             ADDR => address,
               DO => instruction(15 downto 0),
              DOP => instruction(17 downto 16)); 
--
end low_level_definition;
--
------------------------------------------------------------------------------------
--
-- END OF FILE monitor.vhd
--
------------------------------------------------------------------------------------
